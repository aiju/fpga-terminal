library IEEE;
use IEEE.STD_LOGIC_1164.all;

package const is
	constant cols : integer := 80;
	constant lines : integer := 30;
	constant buflines : integer := 50;
end const;

package body const is

end const;
